/*
    CS/ECE 552 FALL '22
    Homework #2, Problem 1

    1 input NOT
*/
module not1 (out, in1);
    output wire out;
    input wire in1;
    assign out = ~in1;
endmodule
